
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity project_tb is
end project_tb;

architecture projecttb of project_tb is
constant c_CLOCK_PERIOD         : time := 15 ns;
signal   tb_done                : std_logic;
signal   mem_address            : std_logic_vector (15 downto 0) := (others => '0');
signal   tb_rst                 : std_logic := '0';
signal   tb_start               : std_logic := '0';
signal   tb_clk                 : std_logic := '0';
signal   mem_o_data,mem_i_data  : std_logic_vector (7 downto 0);
signal   enable_wire            : std_logic;
signal   mem_we                 : std_logic;
signal   i                      : std_logic_vector (1 downto 0)  := std_logic_vector(to_unsigned( 0, 2)); 

type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
signal RAM0: ram_type := (0 => std_logic_vector(to_unsigned( 1, 8)), 
						 1 => std_logic_vector(to_unsigned( 1, 8)), 
						 2 => std_logic_vector(to_unsigned( 0, 8)),
						 others => (others =>'0')); 
signal RAM1: ram_type := (0 => std_logic_vector(to_unsigned( 3, 8)), 
						 1 => std_logic_vector(to_unsigned( 5, 8)), 
						 2 => std_logic_vector(to_unsigned( 1, 8)),
						 3 => std_logic_vector(to_unsigned( 1, 8)),
						 4 => std_logic_vector(to_unsigned( 1, 8)),
						 5 => std_logic_vector(to_unsigned( 0, 8)),
						 6 => std_logic_vector(to_unsigned( 0, 8)),
						 7 => std_logic_vector(to_unsigned( 1, 8)),
						 8 => std_logic_vector(to_unsigned( 0, 8)),
						 9 => std_logic_vector(to_unsigned( 0, 8)),
						 10 => std_logic_vector(to_unsigned( 0, 8)),
						 11 => std_logic_vector(to_unsigned( 0, 8)),
						 12 => std_logic_vector(to_unsigned( 0, 8)),
						 13 => std_logic_vector(to_unsigned( 1, 8)),
						 14 => std_logic_vector(to_unsigned( 1, 8)),
						 15 => std_logic_vector(to_unsigned( 0, 8)),
						 16 => std_logic_vector(to_unsigned( 1, 8)),
						 others => (others =>'0')); 
signal RAM2: ram_type := (0 => std_logic_vector(to_unsigned( 1, 8)), 
						 1 => std_logic_vector(to_unsigned( 1, 8)), 
						 2 => std_logic_vector(to_unsigned( 10, 8)),
						 others => (others =>'0')); 
signal RAM3: ram_type := (0 => std_logic_vector(to_unsigned( 6, 8)), 
						 1 => std_logic_vector(to_unsigned( 2, 8)), 
						 2 => std_logic_vector(to_unsigned( 187, 8)),
						 3 => std_logic_vector(to_unsigned( 233, 8)),
						 4 => std_logic_vector(to_unsigned( 235, 8)),
						 5 => std_logic_vector(to_unsigned( 179, 8)),
						 6 => std_logic_vector(to_unsigned( 166, 8)),
						 7 => std_logic_vector(to_unsigned( 255, 8)),
						 8 => std_logic_vector(to_unsigned( 219, 8)),
						 9 => std_logic_vector(to_unsigned( 0, 8)),
						 10 => std_logic_vector(to_unsigned( 60, 8)),
						 11 => std_logic_vector(to_unsigned( 135, 8)),
						 12 => std_logic_vector(to_unsigned( 12, 8)),
						 13 => std_logic_vector(to_unsigned( 62, 8)),
						 others => (others =>'0')); 

component project_reti_logiche is
port (
      i_clk         : in  std_logic;
      i_start       : in  std_logic;
      i_rst         : in  std_logic;
      i_data        : in  std_logic_vector(7 downto 0);
      o_address     : out std_logic_vector(15 downto 0);
      o_done        : out std_logic;
      o_en          : out std_logic;
      o_we          : out std_logic;
      o_data        : out std_logic_vector (7 downto 0)
      );
end component project_reti_logiche;


begin
UUT: project_reti_logiche
port map (
          i_clk      	=> tb_clk,
          i_start       => tb_start,
          i_rst      	=> tb_rst,
          i_data    	=> mem_o_data,
          o_address  	=> mem_address,
          o_done      	=> tb_done,
          o_en   	    => enable_wire,
          o_we 		    => mem_we,
          o_data    	=> mem_i_data
          );

p_CLK_GEN : process is
begin
    wait for c_CLOCK_PERIOD/2;
    tb_clk <= not tb_clk;
end process p_CLK_GEN;


MEM : process(tb_clk)
begin
	 if tb_clk'event and tb_clk = '1' then
		 if enable_wire = '1' then
			 if i = std_logic_vector(to_unsigned( 0, 2)) then
				 if mem_we = '1' then
					 RAM0(conv_integer(mem_address)) <= mem_i_data;
					 mem_o_data <= mem_i_data after 1 ns;
				 else
					 mem_o_data <= RAM0(conv_integer(mem_address)) after 1 ns;
				 end if;
			 elsif i = std_logic_vector(to_unsigned( 1, 2)) then
				 if mem_we = '1' then
					 RAM1(conv_integer(mem_address)) <= mem_i_data;
					 mem_o_data <= mem_i_data after 1 ns;
				 else
					 mem_o_data <= RAM1(conv_integer(mem_address)) after 1 ns;
				 end if;			 
			 elsif i = std_logic_vector(to_unsigned( 2, 2)) then
				 if mem_we = '1' then
					 RAM2(conv_integer(mem_address)) <= mem_i_data;
					 mem_o_data <= mem_i_data after 1 ns;
				 else
					 mem_o_data <= RAM2(conv_integer(mem_address)) after 1 ns;
				 end if;			 
			 elsif i = std_logic_vector(to_unsigned( 3, 2)) then
				 if mem_we = '1' then
					 RAM3(conv_integer(mem_address)) <= mem_i_data;
					 mem_o_data <= mem_i_data after 1 ns;
				 else
					 mem_o_data <= RAM3(conv_integer(mem_address)) after 1 ns;
				 end if;			 
			 end if;
		 end if;
	 end if;
end process;



test : process is
begin
	 wait for 100 ns;
	 wait for c_CLOCK_PERIOD;
	 tb_rst <= '1';
	 wait for c_CLOCK_PERIOD;
	 wait for 100 ns;
	 tb_rst <= '0';
	 wait for c_CLOCK_PERIOD;
	 wait for 100 ns;
	 tb_start <= '1';
	 wait for c_CLOCK_PERIOD;
	 wait until tb_done = '1';
	 wait for c_CLOCK_PERIOD;
	 tb_start <= '0';
	 wait until tb_done = '0';
	 wait for 100 ns; 
	 
     --
     tb_rst <= '1';
	 wait for c_CLOCK_PERIOD;
	 wait for 100 ns;
	 tb_rst <= '0';
     --
 
     i <= std_logic_vector(to_unsigned( 1, 2));
 	 wait for 100 ns;
	 tb_start <= '1';
	 --
	 wait for 500 ns;
	 tb_rst <= '1';
	 wait for c_CLOCK_PERIOD;
	 wait for 100 ns;
	 tb_rst <= '0';
	 --i <= std_logic_vector(to_unsigned( 2, 2));
	 wait for 100 ns;
	 --
	 
	 wait for c_CLOCK_PERIOD;
	 wait until tb_done = '1';
	 wait for c_CLOCK_PERIOD;
	 tb_start <= '0';
	 wait until tb_done = '0';
	 wait for 100 ns;
	 i <= std_logic_vector(to_unsigned( 3, 2));
 
 	 wait for 100 ns;
	 tb_start <= '1';
	 wait for c_CLOCK_PERIOD;
	 wait until tb_done = '1';
	 wait for c_CLOCK_PERIOD;
	 tb_start <= '0';
	 wait until tb_done = '0';
	 wait for 100 ns;



	 assert RAM0(3) = std_logic_vector(to_unsigned( 0, 8)) report " TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM0(3))))  severity failure; 
  

	 assert RAM2(3) = std_logic_vector(to_unsigned( 0, 8)) report " TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM2(3))))  severity failure; 
 

	 assert RAM3(14) = std_logic_vector(to_unsigned( 187, 8)) report " TEST FALLITO (WORKING ZONE). Expected  187  found " & integer'image(to_integer(unsigned(RAM3(14))))  severity failure; 
 	 assert RAM3(15) = std_logic_vector(to_unsigned( 233, 8)) report " TEST FALLITO (WORKING ZONE). Expected  233  found " & integer'image(to_integer(unsigned(RAM3(15))))  severity failure; 
 	 assert RAM3(16) = std_logic_vector(to_unsigned( 235, 8)) report " TEST FALLITO (WORKING ZONE). Expected  235  found " & integer'image(to_integer(unsigned(RAM3(16))))  severity failure; 
 	 assert RAM3(17) = std_logic_vector(to_unsigned( 179, 8)) report " TEST FALLITO (WORKING ZONE). Expected  179  found " & integer'image(to_integer(unsigned(RAM3(17))))  severity failure; 
 	 assert RAM3(18) = std_logic_vector(to_unsigned( 166, 8)) report " TEST FALLITO (WORKING ZONE). Expected  166  found " & integer'image(to_integer(unsigned(RAM3(18))))  severity failure; 
 	 assert RAM3(19) = std_logic_vector(to_unsigned( 255, 8)) report " TEST FALLITO (WORKING ZONE). Expected  255  found " & integer'image(to_integer(unsigned(RAM3(19))))  severity failure; 
 	 assert RAM3(20) = std_logic_vector(to_unsigned( 219, 8)) report " TEST FALLITO (WORKING ZONE). Expected  219  found " & integer'image(to_integer(unsigned(RAM3(20))))  severity failure; 
 	 assert RAM3(21) = std_logic_vector(to_unsigned( 0, 8)) report " TEST FALLITO (WORKING ZONE). Expected  0  found " & integer'image(to_integer(unsigned(RAM3(21))))  severity failure; 
 	 assert RAM3(22) = std_logic_vector(to_unsigned( 60, 8)) report " TEST FALLITO (WORKING ZONE). Expected  60  found " & integer'image(to_integer(unsigned(RAM3(22))))  severity failure; 
 	 assert RAM3(23) = std_logic_vector(to_unsigned( 135, 8)) report " TEST FALLITO (WORKING ZONE). Expected  135  found " & integer'image(to_integer(unsigned(RAM3(23))))  severity failure; 
 	 assert RAM3(24) = std_logic_vector(to_unsigned( 12, 8)) report " TEST FALLITO (WORKING ZONE). Expected  12  found " & integer'image(to_integer(unsigned(RAM3(24))))  severity failure; 
 	 assert RAM3(25) = std_logic_vector(to_unsigned( 62, 8)) report " TEST FALLITO (WORKING ZONE). Expected  62  found " & integer'image(to_integer(unsigned(RAM3(25))))  severity failure; 
 

    assert false report "Simulation Ended! TEST PASSATO" severity failure;
end process test;

end projecttb; 